`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    20:06:47 01/02/2017 
// Design Name: 
// Module Name:    cars 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module cars(
    output wire red_car1,
    output wire red_car2,
    output wire yellow_car1,
    output wire yellow_car2, 
	output wire signed [11:0]car1_s,
	output wire signed [11:0]car1_e,
	output wire signed [11:0]car2_s,
	output wire signed [11:0]car2_e,
	output wire signed [11:0]car3_s,
	output wire signed [11:0]car3_e,
	output wire signed [11:0]car4_s,
	output wire signed [11:0]car4_e,
	input clk,
  	input rst,
    input [23:0]sec_count,
    input [10:0]col,
    input [10:0]row
    );




wire [159:0]red_car[0:59];

assign red_car[0]  = 160'b0000001111111111111111111111111111111111000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000;
assign red_car[1]  = 160'b0000111111111111111111111111111111111110001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000;
assign red_car[2]  = 160'b0011111111111111111111111111111111111100011100000011111111100000011111111100000000000111111111111111111111111111111111111111111111111111111111111111111111111100;
assign red_car[3]  = 160'b0011111111111111111111111111111111111000100000000001111000000111000011110000001111000001111111111111111111111111111111111111111111111111111111111111111111111100;
assign red_car[4]  = 160'b0111111111111111111111111111111111110000000011111000000001111111111000000001111111111000000000111111111111111111111111111111111111111111111111111111111111111110;
assign red_car[5]  = 160'b0111111111111111111111111111111111100001111111111111111111111111111111111111111111111111100000000011111111111111111111111111111111111111111111111111111111111110;
assign red_car[6]  = 160'b1111111111111111111111111111111111000001111111111111111111111111111111111111111111111111111100000000111111111111111111111111111111111111111111111111111111111111;
assign red_car[7]  = 160'b1111111111111111111111111111111111000011111111111111111111111111111111111111111111111111111111111000000001111111111111111111111111111111111111111111111111111111;
assign red_car[8]  = 160'b1111111111111111111111111111111110000011111111111111111111111111111111111111111111111111111111111111100000000111111111111111111111111111111111111111111111111111;
assign red_car[9]  = 160'b1111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
assign red_car[10] = 160'b1111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
assign red_car[11] = 160'b1111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
assign red_car[12] = 160'b1111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
assign red_car[13] = 160'b1111111111111111111111111111110000001111111111111111110000000111111111111111111111111111111111111111111111111111111111111111111111000000000000111111111111111111;
assign red_car[14] = 160'b0011111111111111111111111111110000011111111111111111111111000000000011111111111111111111111111111111111111111111111111111111110000000000000111111111111111111111;
assign red_car[15] = 160'b0000111111111111111111111111100000011111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111;
assign red_car[16] = 160'b0000011111111111111111111111100000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
assign red_car[17] = 160'b0000001111111111111111111111000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
assign red_car[18] = 160'b0000001111111111111111111111000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
assign red_car[19] = 160'b0000001111111111111111111110000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
assign red_car[20] = 160'b0000001111111111111111111110000000111111111110000000000111111111111111111111100000111111111111111000000001111111111111111111000000011111111111111111111111111111;
assign red_car[21] = 160'b0000001111111111111111111110000000111111110000000000000111111111111111111110000000011111111111111000000001111111111111110000000000011111111111111111111111111111;
assign red_car[22] = 160'b0000011111111111111111111100000000111111000011111110000111111111111111111100011110001111111111111000000001111111111111000011111000011111111111111111111111111111;
assign red_car[23] = 160'b0000111111111111111111111100000000111100000011111111000111111111111111111000111111000111111111111000000001111111111100000111111000011111111111111111111111111111;
assign red_car[24] = 160'b0011111111111111111111111100000000111111000011111111000111111111111111110001111111100011111111111000000001111111111100001111111000011111111111111111111111111111;
assign red_car[25] = 160'b1111111111111111111111111100000000111111100000000000000111111111111111100000000000000001111111111000000001111111111100001111111000011111111111111111111111111111;
assign red_car[26] = 160'b1111111111111111111111111100000000111111100000000001000111111111111111000000000000000000111111111000000001111111111110000111111000011111111111111111111111111111;
assign red_car[27] = 160'b1111111111111111111111111100000000111111000011111111000111111111111110001111111111111100011111111000000001111111111110000011111000011111111111111111111111111111;
assign red_car[28] = 160'b1111111111111111111111111100000000111100000111111111000111111111111100011111111111111110001111111000000001111111111111100000111000011111111111111111111111111111;
assign red_car[29] = 160'b1111111111111111111111111100000000111000000111111111000111111111111000111111111111111111000111111000000001111111111111111100000000011111111111111111111111111111;
assign red_car[30] = 160'b1111111111111111111111111100000000111110000000000001000111111111110001111111111111111111100011111000000001111111111111111111100000011111111111111111111111111111;
assign red_car[31] = 160'b1111111111111111111111111100000000111111111111111111111111111111111111111111111111111111111111111000000001111111111111111111111111111111111111111111111111111111;
assign red_car[32] = 160'b1111111111111111111111111100000000111111111111111111111111111111111111111111111111111111111111111000000001111111111111111111111111111111111111111111111111111111;
assign red_car[33] = 160'b1111111111111111111111111100000000111111111111111111111111111111111111111111111111111111111111111000000001111111111111111111111111111111111111111111111111111111;
assign red_car[34] = 160'b1111111111111111111111111100000000111111111111111111111111111111111111111111111111111111111111111000000001111111111111111111111111111111111111111111111111111111;
assign red_car[35] = 160'b0011111111111111111111111100000000111111111111111111000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111;
assign red_car[36] = 160'b0000111111111111111111111100000000111111111111111111000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111;
assign red_car[37] = 160'b0000011111111111111111111100000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
assign red_car[38] = 160'b0000001111111111111111111110000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
assign red_car[39] = 160'b0000001111111111111111111110000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
assign red_car[40] = 160'b0000001111111111111111111110000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
assign red_car[41] = 160'b0000001111111111111111111111000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
assign red_car[42] = 160'b0000001111111111111111111111000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
assign red_car[43] = 160'b0000011111111111111111111111100000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
assign red_car[44] = 160'b0000111111111111111111111111100000011111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111;
assign red_car[45] = 160'b0011111111111111111111111111110000011111111111111111111111000000000011111111111111111111111111111111111111111111111111111111110000000000000111111111111111111111;
assign red_car[46] = 160'b1111111111111111111111111111110000001111111111111111110000000111111111111111111111111111111111111111111111111111111111111111111111000000000000111111111111111111;
assign red_car[47] = 160'b1111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
assign red_car[48] = 160'b1111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
assign red_car[49] = 160'b1111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
assign red_car[50] = 160'b1111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
assign red_car[51] = 160'b1111111111111111111111111111111110000011111111111111111111111111111111111111111111111111111111111111100000000111111111111111111111111111111111111111111111111111;
assign red_car[52] = 160'b1111111111111111111111111111111111000011111111111111111111111111111111111111111111111111111111111000000001111111111111111111111111111111111111111111111111111111;
assign red_car[53] = 160'b1111111111111111111111111111111111000001111111111111111111111111111111111111111111111111111100000000111111111111111111111111111111111111111111111111111111111111;
assign red_car[54] = 160'b0111111111111111111111111111111111100001111111111111111111111111111111111111111111111111100000000011111111111111111111111111111111111111111111111111111111111110;
assign red_car[55] = 160'b0111111111111111111111111111111111110000000011111000000001111111111000000001111111111000000000111111111111111111111111111111111111111111111111111111111111111110;
assign red_car[56] = 160'b0011111111111111111111111111111111111000100000000001111000000111000011110000001111000001111111111111111111111111111111111111111111111111111111111111111111111100;
assign red_car[57] = 160'b0011111111111111111111111111111111111100011100000011111111100000011111111100000000000111111111111111111111111111111111111111111111111111111111111111111111111100;
assign red_car[58] = 160'b0000111111111111111111111111111111111110001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000;
assign red_car[59] = 160'b0000001111111111111111111111111111111111000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000;




reg [5:0]red_car_count;
reg [159:0]red_car_pix;

reg signed[11:0]red_car_flag1;
reg signed[11:0]red_car_start1;
reg signed[11:0]red_car_end1;

reg signed[11:0]red_car_flag2;
reg signed[11:0]red_car_start2;
reg signed[11:0]red_car_end2;


always@(posedge clk or posedge rst)
  if(rst)                                          red_car_count<=0;
  else if(row>510)                             red_car_count<=0;
  else if(row>450 && row <=510 && col==1000) red_car_count<=red_car_count+1;
  else                                             red_car_count<=red_car_count;
  
always@(posedge clk or posedge rst)
  if(rst)                                          red_car_pix<=0;
  else if(row>450 && row <=510)             red_car_pix<=red_car[red_car_count];
  else                                             red_car_pix<=0;    

always@(posedge clk or posedge rst)
  if(rst) red_car_flag1=0;
  else if(sec_count==0)
    if(red_car_flag1<=180) red_car_flag1=red_car_flag1+6;
    else red_car_flag1 = -779;
  else red_car_flag1=red_car_flag1;
  
always@(posedge clk or posedge rst)
  if(rst) red_car_flag2=0;
  else if(sec_count==0)
    if(red_car_flag2<=580) red_car_flag2=red_car_flag2+6;
    else red_car_flag2 = -379;
  else red_car_flag2=red_car_flag2;




always@(posedge clk or posedge rst)
  if(rst) begin
    red_car_start1=620;
    red_car_end1=779;
  end
  else begin
    red_car_start1=620+red_car_flag1;
    red_car_end1=779+red_car_flag1;
  end
  
always@(posedge clk or posedge rst)
  if(rst) begin
    red_car_start2=220;
    red_car_end2=379;
  end
  else begin
    red_car_start2=220+red_car_flag2;
    red_car_end2=379+red_car_flag2;
  end
  
wire signed[11:0]temp1;
wire signed[11:0]temp2;


assign temp1=(red_car_start1<=0)?0:red_car_start1;
assign temp2=(red_car_start2<=0)?0:red_car_start2;


assign red_car1=(row>450 && row <=510 && temp1+104<=col && red_car_end1+104 >=col)?red_car_pix[col-red_car_end1-104+159]:0;
assign red_car2=(row>450 && row <=510 && temp2+104<=col && red_car_end2+104 >=col)?red_car_pix[col-red_car_end2-104+159]:0;



reg [5:0]yellow_car_count;
reg [0:159]yellow_car_pix;



reg signed[11:0]yellow_car_flag1;
reg signed[11:0]yellow_car_start1;
reg signed[11:0]yellow_car_end1;

reg signed[11:0]yellow_car_flag2;
reg signed[11:0]yellow_car_start2;
reg signed[11:0]yellow_car_end2;

assign car1_s=red_car_start1+104;
assign car1_e=red_car_end1+104;
assign car2_s=red_car_start2+104;
assign car2_e=red_car_end2+104;
assign car3_s=yellow_car_start1+104;
assign car3_e=yellow_car_end1+104;
assign car4_s=yellow_car_start2+104;
assign car4_e=yellow_car_end2+104;

always@(posedge clk or posedge rst)
  if(rst)                                          yellow_car_count<=0;
  else if(row>430)                             yellow_car_count<=0;
  else if(row>370 && row <=430 && col==1000) yellow_car_count<=yellow_car_count+1;
  else                                             yellow_car_count<=yellow_car_count;

always@(posedge clk or posedge rst)
  if(rst)                                          yellow_car_pix<=0;
  else if(row>370 && row <=430)             yellow_car_pix<=red_car[yellow_car_count];
  else                                             yellow_car_pix<=0;    

always@(posedge clk or posedge rst)
  if(rst)                       yellow_car_flag1=0;
  else if(sec_count==0)
      if(yellow_car_flag1>=-459)yellow_car_flag1=yellow_car_flag1-8;
      else                      yellow_car_flag1 = 500;
  else                          yellow_car_flag1=yellow_car_flag1;
  
always@(posedge clk or posedge rst)
  if(rst)                       yellow_car_flag2=0;
  else if(sec_count==0)
    if(yellow_car_flag2>=-779)  yellow_car_flag2=yellow_car_flag2-8;
    else                        yellow_car_flag2 = 180;
  else                          yellow_car_flag2=yellow_car_flag2;



always@(posedge clk or posedge rst)
  if(rst) begin
    yellow_car_start1=300;
    yellow_car_end1=459;
  end
  else begin
    yellow_car_start1=300+yellow_car_flag1;
    yellow_car_end1=459+yellow_car_flag1;
  end
  
always@(posedge clk or posedge rst)
  if(rst) begin
    yellow_car_start2=620;
    yellow_car_end2=779;
  end
  else begin
    yellow_car_start2=620+yellow_car_flag2;
    yellow_car_end2=779+yellow_car_flag2;
  end
  
wire signed[11:0]temp3;
wire signed[11:0]temp4;


assign temp3=(yellow_car_end1>=800)?800:yellow_car_end1;
assign temp4=(yellow_car_end2>=800)?800:yellow_car_end2;


assign yellow_car1=(row>370 && row <=430 && yellow_car_start1+104<=col && temp3+104 >=col)?yellow_car_pix[col-yellow_car_end1-104+159]:0;
assign yellow_car2=(row>370 && row <=430 && yellow_car_start2+104<=col && temp4+104 >=col)?yellow_car_pix[col-yellow_car_end2-104+159]:0;



endmodule
